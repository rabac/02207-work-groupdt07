entity and_or_inv is
  port ( a1, a2, b1, b2 : in bit := '1';
	 y : out bit );
end entity and_or_inv;
