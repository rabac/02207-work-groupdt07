entity ap_a_10 is

end entity ap_a_10;


library ieee;  use ieee.std_logic_1164.all;
library util;  use util.stimulus_generators.all;

architecture test of ap_a_10 is

  signal a, b, c, d : std_ulogic;
  signal test_vector : std_ulogic_vector(1 to 4);

begin

  b1 : block is
    signal y : std_ulogic;
  begin
    -- code from book

    y <= a or b or c or d;

    -- end code from book
  end block b1;

  b2 : block is
    signal y : std_ulogic;
  begin
    -- code from book

    y <= ( a or b ) or ( c or d );

    -- end code from book
  end block b2;

  b3 : block is
    signal y : std_ulogic;
  begin
    -- code from book (syntax error)

    -- y <= a or b or c and d;

    -- end code from book
  end block b3;

  b4 : block is
    signal y : std_ulogic;
  begin
    -- code from book

    y <= ( a or b ) or ( c and d );

    -- end code from book
  end block b4;

  stimulus : all_possible_values(test_vector, 10 ns);

  (a, b, c, d) <= test_vector;

end architecture test;

