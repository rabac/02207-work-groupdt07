package ch_05_19 is

  -- code from book:

  subtype digit is bit_vector(3 downto 0);

  -- end of code from book

end package ch_05_19;
