entity fg_a_01 is
end entity fg_a_01;



library ieee;  use ieee.std_logic_1164.all;

architecture test of fg_a_01 is

  signal clk, d : std_ulogic;

begin

  stimulus : process is
  begin
    clk <= '0';  d <= '0';  wait for 10 ns;
    clk <= '1', '0' after 10 ns;  wait for 20 ns;
    d <= '1';  wait for 10 ns;
    clk <= '1', '0' after 20 ns;  d <= '0' after 10 ns;

    wait;
  end process stimulus;


  b1 : block is
    signal q : std_ulogic;
  begin

  -- code from book

process (clk) is
begin
  if rising_edge(clk) then
    q <= d;
  end if;
end process;

  -- end code from book

  end block b1;


  b2 : block is
    signal q : std_ulogic;
  begin

  -- code from book

process is
begin
  wait until rising_edge(clk);
  q <= d;
end process;

  -- end code from book

  end block b2;


  b3 : block is
    signal q : std_ulogic;
  begin

  -- code from book

q <= d when rising_edge(clk) else
    q;

  -- end code from book

  end block b3;


  b4 : block is
    signal q : std_ulogic;
  begin

  -- code from book

b : block ( rising_edge(clk)
            and not clk'stable ) is
begin
  q <= guarded d;
end block b;

  -- end code from book

  end block b4;

end architecture test;
