entity ap_a_06 is

end entity ap_a_06;


library ieee;  use ieee.std_logic_1164.all;

architecture test of ap_a_06 is

  signal a, ts, x : std_ulogic;

begin

  -- code from book

  ts <= a when x = '1' else
        'Z';

  -- end code from book

  x <= '0', '1' after 20 ns;
  a <= '0', '1' after 10 ns, '0' after 20 ns, '1' after 30 ns;

end architecture test;

