entity to_vector_test is

end entity to_vector_test;
