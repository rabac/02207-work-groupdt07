library ieee;  use ieee.std_logic_1164.all;

package alu_types is

  subtype alu_func is std_ulogic_vector(3 downto 0);

  constant alu_add : alu_func := "0000";
  constant alu_addu : alu_func := "0001";
  constant alu_sub : alu_func := "0010";
  constant alu_subu : alu_func := "0011";

end package alu_types;
