entity fg_a_06 is

end entity fg_a_06;


library ieee;  use ieee.std_logic_1164.all;

architecture test of fg_a_06 is

  -- code from book

  constant terminal_count : integer := 2**6 - 1;
  subtype counter_range is integer range 0 to terminal_count;
  signal count : counter_range;
  -- . . .

  -- end code from book

  signal clk, reset : std_ulogic;

begin

  -- code from book

  counter6 : process (reset, clk)
  begin
    if reset = '0' then
      count <= 0;
    elsif rising_edge(clk) then
      if count < terminal_count then
        count <= count + 1;
      else
        count <= 0;
      end if;
    end if;
  end process counter6;

  -- end code from book

  stimulus : process is
  begin
    reset <= '1';  clk <= '0';  wait for 10 ns;
    clk <= '1', '0' after 10 ns;  wait for 20 ns;
    clk <= '1', '0' after 10 ns;  wait for 20 ns;
    clk <= '1', '0' after 10 ns;  wait for 20 ns;
    reset <= '0', '1' after 30 ns;
    clk <= '1' after 10 ns, '0' after 20 ns;
    wait for 40 ns;
    for i in 1 to terminal_count + 10 loop
      clk <= '1', '0' after 10 ns;
      wait for 20 ns;
    end loop;

    wait;
  end process stimulus;

end architecture test;

