entity fg_a_04 is

end entity fg_a_04;


library ieee;  use ieee.std_logic_1164.all;

architecture test of fg_a_04 is

  signal clk, reset, d, q, q_n : std_ulogic;

begin

  -- code from book

  ff1 : process (reset, clk) is
  begin
    if reset = '1' then
      q <= '0';
    elsif rising_edge(clk) then
      q <= d;
    end if;
  end process ff1;

  q_n <= not q;

  -- end code from book

  stimulus : process is
  begin
    reset <= '0';  clk <= '0';  d <= '1';  wait for 10 ns;
    reset <= '1', '0' after 30 ns;
    clk <= '1' after 10 ns, '0' after 20 ns;
    wait for 40 ns;
    clk <= '1', '0' after 20 ns;
    d <= '0' after 10 ns;

    wait;
  end process stimulus;

end architecture test;

