entity dlx_test is

end entity dlx_test;
