library ieee;  use ieee.std_logic_1164.std_ulogic;

entity logic_block is
  port ( a, b : in std_ulogic;
         y, z : out std_ulogic );
end entity logic_block;
