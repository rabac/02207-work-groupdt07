entity bv_test is
  
end entity bv_test;
