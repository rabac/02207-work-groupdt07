-- not in book

use work.tb_05_13.all;

-- end not in book

entity adder is
  port ( a, b : in word;
         sum : out word );
end entity adder;
