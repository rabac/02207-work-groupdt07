package tb_05_13 is

  subtype word is integer;

end package tb_05_13;
