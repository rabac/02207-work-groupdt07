entity test_bench_04_03 is

end entity test_bench_04_03;


----------------------------------------------------------------


use work.pk_04_02.all;


architecture test_byte_swap_behavior of test_bench_04_03 is

  signal input, output : halfword := x"0000";

begin

  dut : entity work.byte_swap(behavior)
    port map ( input => input, output => output );

  stumulus : process is
  begin
			wait for 10 ns;
    input <= x"ff00";	wait for 10 ns;
    input <= x"00ff";	wait for 10 ns;
    input <= x"aa33";	wait for 10 ns;

    wait;
  end process stumulus;

end architecture test_byte_swap_behavior;
