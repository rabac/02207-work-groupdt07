entity multiplier_test is

end entity multiplier_test;
