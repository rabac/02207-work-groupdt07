entity ent is

end entity ent;
