entity ap_a_01 is

end entity ap_a_01;


library ieee;  use ieee.std_logic_1164.all;

architecture test of ap_a_01 is

  signal clk : std_ulogic;

begin

  process (clk) is

    -- code from book

    -- end code from book

  begin

    if

    -- code from book

    clk'event and (To_X01(clk) = '1') and (To_X01(clk'last_value) = '0')

    -- end code from book

    then
      report "rising edge on clk";
    end if;

  end process;

  clk <= '0', '1' after 10 ns, '0' after 20 ns,
         '1' after 30 ns, '0' after 40 ns;

end architecture test;

