entity ap_a_05 is

end entity ap_a_05;


library ieee;  use ieee.std_logic_1164.all;

architecture test of ap_a_05 is

  signal a, b, y, x : std_ulogic;

begin

  -- code from book

  y <= a when x = '1' else
       b;

  -- end code from book

  x <= '0', '1' after 20 ns;
  a <= '0', '1' after 10 ns, '0' after 20 ns, '1' after 30 ns;
  b <= '0', '1' after 15 ns, '0' after 25 ns, '1' after 35 ns;

end architecture test;

